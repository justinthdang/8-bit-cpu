library verilog;
use verilog.vl_types.all;
entity ssegreport_vlg_vec_tst is
end ssegreport_vlg_vec_tst;
