library verilog;
use verilog.vl_types.all;
entity regreport_vlg_vec_tst is
end regreport_vlg_vec_tst;
