library verilog;
use verilog.vl_types.all;
entity fsmreport_vlg_vec_tst is
end fsmreport_vlg_vec_tst;
