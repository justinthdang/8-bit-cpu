library verilog;
use verilog.vl_types.all;
entity test3_vlg_vec_tst is
end test3_vlg_vec_tst;
