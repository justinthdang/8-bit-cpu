library verilog;
use verilog.vl_types.all;
entity dec3to8report_vlg_vec_tst is
end dec3to8report_vlg_vec_tst;
